module Register_Bunch(
    input   
);