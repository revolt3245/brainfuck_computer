module ALU(

);

endmodule;